module mu0 (
    input clk
);

endmodule
